magic
tech sky130A
magscale 1 2
timestamp 1729701459
<< obsli1 >>
rect 13104 5159 570808 352809
<< obsm1 >>
rect 13104 8 570808 352840
<< metal2 >>
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
<< obsm2 >>
rect 386 536 577382 352829
rect 386 2 486 536
rect 710 2 1590 536
rect 1814 2 125790 536
rect 126014 2 126894 536
rect 127118 2 129286 536
rect 129510 2 130482 536
rect 130706 2 132874 536
rect 133098 2 134070 536
rect 134294 2 136370 536
rect 136594 2 137566 536
rect 137790 2 139958 536
rect 140182 2 141154 536
rect 141378 2 143454 536
rect 143678 2 144650 536
rect 144874 2 147042 536
rect 147266 2 148238 536
rect 148462 2 150538 536
rect 150762 2 151734 536
rect 151958 2 154126 536
rect 154350 2 155322 536
rect 155546 2 157714 536
rect 157938 2 158818 536
rect 159042 2 161210 536
rect 161434 2 162406 536
rect 162630 2 164798 536
rect 165022 2 165994 536
rect 166218 2 168294 536
rect 168518 2 169490 536
rect 169714 2 171882 536
rect 172106 2 173078 536
rect 173302 2 175378 536
rect 175602 2 176574 536
rect 176798 2 178966 536
rect 179190 2 180162 536
rect 180386 2 182462 536
rect 182686 2 183658 536
rect 183882 2 186050 536
rect 186274 2 187246 536
rect 187470 2 189638 536
rect 189862 2 190742 536
rect 190966 2 193134 536
rect 193358 2 194330 536
rect 194554 2 196722 536
rect 196946 2 197826 536
rect 198050 2 200218 536
rect 200442 2 201414 536
rect 201638 2 203806 536
rect 204030 2 205002 536
rect 205226 2 207302 536
rect 207526 2 208498 536
rect 208722 2 210890 536
rect 211114 2 212086 536
rect 212310 2 214386 536
rect 214610 2 215582 536
rect 215806 2 217974 536
rect 218198 2 219170 536
rect 219394 2 221470 536
rect 221694 2 222666 536
rect 222890 2 225058 536
rect 225282 2 226254 536
rect 226478 2 228646 536
rect 228870 2 229750 536
rect 229974 2 232142 536
rect 232366 2 233338 536
rect 233562 2 235730 536
rect 235954 2 236926 536
rect 237150 2 239226 536
rect 239450 2 240422 536
rect 240646 2 242814 536
rect 243038 2 244010 536
rect 244234 2 246310 536
rect 246534 2 247506 536
rect 247730 2 249898 536
rect 250122 2 251094 536
rect 251318 2 253394 536
rect 253618 2 254590 536
rect 254814 2 256982 536
rect 257206 2 258178 536
rect 258402 2 260570 536
rect 260794 2 261674 536
rect 261898 2 264066 536
rect 264290 2 265262 536
rect 265486 2 267654 536
rect 267878 2 268758 536
rect 268982 2 271150 536
rect 271374 2 272346 536
rect 272570 2 274738 536
rect 274962 2 275934 536
rect 276158 2 278234 536
rect 278458 2 279430 536
rect 279654 2 281822 536
rect 282046 2 283018 536
rect 283242 2 285318 536
rect 285542 2 286514 536
rect 286738 2 288906 536
rect 289130 2 290102 536
rect 290326 2 292494 536
rect 292718 2 293598 536
rect 293822 2 295990 536
rect 296214 2 297186 536
rect 297410 2 299578 536
rect 299802 2 300682 536
rect 300906 2 303074 536
rect 303298 2 304270 536
rect 304494 2 306662 536
rect 306886 2 307858 536
rect 308082 2 310158 536
rect 310382 2 311354 536
rect 311578 2 313746 536
rect 313970 2 314942 536
rect 315166 2 317242 536
rect 317466 2 318438 536
rect 318662 2 320830 536
rect 321054 2 322026 536
rect 322250 2 324326 536
rect 324550 2 325522 536
rect 325746 2 327914 536
rect 328138 2 329110 536
rect 329334 2 331502 536
rect 331726 2 332606 536
rect 332830 2 334998 536
rect 335222 2 336194 536
rect 336418 2 338586 536
rect 338810 2 339782 536
rect 340006 2 342082 536
rect 342306 2 343278 536
rect 343502 2 345670 536
rect 345894 2 346866 536
rect 347090 2 349166 536
rect 349390 2 350362 536
rect 350586 2 352754 536
rect 352978 2 353950 536
rect 354174 2 356250 536
rect 356474 2 357446 536
rect 357670 2 359838 536
rect 360062 2 361034 536
rect 361258 2 363426 536
rect 363650 2 364530 536
rect 364754 2 366922 536
rect 367146 2 368118 536
rect 368342 2 370510 536
rect 370734 2 371614 536
rect 371838 2 374006 536
rect 374230 2 375202 536
rect 375426 2 377594 536
rect 377818 2 378790 536
rect 379014 2 381090 536
rect 381314 2 382286 536
rect 382510 2 384678 536
rect 384902 2 385874 536
rect 386098 2 388174 536
rect 388398 2 389370 536
rect 389594 2 391762 536
rect 391986 2 392958 536
rect 393182 2 395258 536
rect 395482 2 396454 536
rect 396678 2 398846 536
rect 399070 2 400042 536
rect 400266 2 402434 536
rect 402658 2 403538 536
rect 403762 2 405930 536
rect 406154 2 407126 536
rect 407350 2 409518 536
rect 409742 2 410714 536
rect 410938 2 413014 536
rect 413238 2 414210 536
rect 414434 2 416602 536
rect 416826 2 417798 536
rect 418022 2 420098 536
rect 420322 2 421294 536
rect 421518 2 423686 536
rect 423910 2 424882 536
rect 425106 2 427182 536
rect 427406 2 428378 536
rect 428602 2 430770 536
rect 430994 2 431966 536
rect 432190 2 434358 536
rect 434582 2 435462 536
rect 435686 2 437854 536
rect 438078 2 439050 536
rect 439274 2 441442 536
rect 441666 2 442546 536
rect 442770 2 444938 536
rect 445162 2 446134 536
rect 446358 2 448526 536
rect 448750 2 449722 536
rect 449946 2 452022 536
rect 452246 2 453218 536
rect 453442 2 455610 536
rect 455834 2 456806 536
rect 457030 2 459106 536
rect 459330 2 460302 536
rect 460526 2 462694 536
rect 462918 2 463890 536
rect 464114 2 466190 536
rect 466414 2 467386 536
rect 467610 2 469778 536
rect 470002 2 470974 536
rect 471198 2 473366 536
rect 473590 2 474470 536
rect 474694 2 476862 536
rect 477086 2 478058 536
rect 478282 2 480450 536
rect 480674 2 481646 536
rect 481870 2 483946 536
rect 484170 2 485142 536
rect 485366 2 487534 536
rect 487758 2 488730 536
rect 488954 2 491030 536
rect 491254 2 492226 536
rect 492450 2 494618 536
rect 494842 2 495814 536
rect 496038 2 498114 536
rect 498338 2 499310 536
rect 499534 2 501702 536
rect 501926 2 502898 536
rect 503122 2 505290 536
rect 505514 2 506394 536
rect 506618 2 508786 536
rect 509010 2 509982 536
rect 510206 2 512374 536
rect 512598 2 513478 536
rect 513702 2 515870 536
rect 516094 2 517066 536
rect 517290 2 519458 536
rect 519682 2 520654 536
rect 520878 2 522954 536
rect 523178 2 524150 536
rect 524374 2 526542 536
rect 526766 2 527738 536
rect 527962 2 530038 536
rect 530262 2 531234 536
rect 531458 2 533626 536
rect 533850 2 534822 536
rect 535046 2 537122 536
rect 537346 2 538318 536
rect 538542 2 540710 536
rect 540934 2 541906 536
rect 542130 2 544298 536
rect 544522 2 545402 536
rect 545626 2 547794 536
rect 548018 2 548990 536
rect 549214 2 551382 536
rect 551606 2 552578 536
rect 552802 2 554878 536
rect 555102 2 556074 536
rect 556298 2 558466 536
rect 558690 2 559662 536
rect 559886 2 561962 536
rect 562186 2 563158 536
rect 563382 2 565550 536
rect 565774 2 566746 536
rect 566970 2 569046 536
rect 569270 2 570242 536
rect 570466 2 572634 536
rect 572858 2 573830 536
rect 574054 2 576222 536
rect 576446 2 577326 536
<< obsm3 >>
rect 381 35 577195 352825
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -7654 2414 711590
rect 5514 -7654 6134 711590
rect 9234 -7654 9854 711590
rect 12954 -7654 13574 711590
rect 16674 -7654 17294 711590
rect 20394 -7654 21014 711590
rect 24114 -7654 24734 711590
rect 27834 -7654 28454 711590
rect 37794 -7654 38414 711590
rect 41514 -7654 42134 711590
rect 45234 -7654 45854 711590
rect 48954 -7654 49574 711590
rect 52674 -7654 53294 711590
rect 56394 -7654 57014 711590
rect 60114 -7654 60734 711590
rect 63834 -7654 64454 711590
rect 73794 -7654 74414 711590
rect 77514 354980 78134 711590
rect 81234 -7654 81854 711590
rect 84954 -7654 85574 711590
rect 88674 -7654 89294 711590
rect 92394 354980 93014 711590
rect 96114 -7654 96734 711590
rect 99834 -7654 100454 711590
rect 109794 -7654 110414 711590
rect 113514 -7654 114134 711590
rect 117234 -7654 117854 711590
rect 120954 -7654 121574 711590
rect 124674 -7654 125294 711590
rect 128394 -7654 129014 711590
rect 132114 -7654 132734 711590
rect 135834 -7654 136454 711590
rect 145794 -7654 146414 711590
rect 149514 -7654 150134 711590
rect 153234 -7654 153854 711590
rect 156954 -7654 157574 711590
rect 160674 -7654 161294 711590
rect 164394 -7654 165014 711590
rect 168114 -7654 168734 711590
rect 171834 -7654 172454 711590
rect 181794 -7654 182414 711590
rect 185514 354980 186134 711590
rect 189234 -7654 189854 711590
rect 192954 -7654 193574 711590
rect 196674 -7654 197294 711590
rect 200394 354980 201014 711590
rect 204114 -7654 204734 711590
rect 207834 -7654 208454 711590
rect 217794 -7654 218414 711590
rect 221514 -7654 222134 711590
rect 225234 -7654 225854 711590
rect 228954 -7654 229574 711590
rect 232674 -7654 233294 711590
rect 236394 -7654 237014 711590
rect 240114 -7654 240734 711590
rect 243834 -7654 244454 711590
rect 253794 -7654 254414 711590
rect 257514 -7654 258134 711590
rect 261234 354980 261854 711590
rect 264954 -7654 265574 711590
rect 268674 -7654 269294 711590
rect 272394 -7654 273014 711590
rect 276114 -7654 276734 711590
rect 279834 -7654 280454 711590
rect 289794 -7654 290414 711590
rect 293514 -7654 294134 711590
rect 297234 -7654 297854 711590
rect 300954 -7654 301574 711590
rect 304674 -7654 305294 711590
rect 308394 354980 309014 711590
rect 312114 -7654 312734 711590
rect 315834 -7654 316454 711590
rect 325794 -7654 326414 711590
rect 329514 -7654 330134 711590
rect 333234 -7654 333854 711590
rect 336954 -7654 337574 711590
rect 340674 -7654 341294 711590
rect 344394 -7654 345014 711590
rect 348114 -7654 348734 711590
rect 351834 -7654 352454 711590
rect 361794 -7654 362414 711590
rect 365514 -7654 366134 711590
rect 369234 354980 369854 711590
rect 372954 -7654 373574 711590
rect 376674 -7654 377294 711590
rect 380394 -7654 381014 711590
rect 384114 354980 384734 711590
rect 387834 -7654 388454 711590
rect 397794 -7654 398414 711590
rect 401514 -7654 402134 711590
rect 405234 -7654 405854 711590
rect 408954 -7654 409574 711590
rect 412674 -7654 413294 711590
rect 416394 -7654 417014 711590
rect 420114 -7654 420734 711590
rect 423834 -7654 424454 711590
rect 433794 -7654 434414 711590
rect 437514 -7654 438134 711590
rect 441234 -7654 441854 711590
rect 444954 -7654 445574 711590
rect 448674 -7654 449294 711590
rect 452394 -7654 453014 711590
rect 456114 -7654 456734 711590
rect 459834 -7654 460454 711590
rect 469794 -7654 470414 711590
rect 473514 -7654 474134 711590
rect 477234 354980 477854 711590
rect 480954 -7654 481574 711590
rect 484674 -7654 485294 711590
rect 488394 -7654 489014 711590
rect 492114 354980 492734 711590
rect 495834 -7654 496454 711590
rect 505794 -7654 506414 711590
rect 509514 -7654 510134 711590
rect 513234 -7654 513854 711590
rect 516954 -7654 517574 711590
rect 520674 -7654 521294 711590
rect 524394 -7654 525014 711590
rect 528114 -7654 528734 711590
rect 531834 -7654 532454 711590
rect 541794 -7654 542414 711590
rect 545514 -7654 546134 711590
rect 549234 -7654 549854 711590
rect 552954 -7654 553574 711590
rect 556674 -7654 557294 711590
rect 560394 -7654 561014 711590
rect 564114 -7654 564734 711590
rect 567834 -7654 568454 711590
rect 577794 -7654 578414 711590
rect 581514 -7654 582134 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 16208 5128 16594 352840
rect 17374 5128 20314 352840
rect 21094 5128 24034 352840
rect 24814 5128 27754 352840
rect 28534 5128 37714 352840
rect 38494 5128 41434 352840
rect 42214 5128 45154 352840
rect 45934 5128 48874 352840
rect 49654 5128 52594 352840
rect 53374 5128 56314 352840
rect 57094 5128 60034 352840
rect 60814 5128 63754 352840
rect 64534 5128 73714 352840
rect 74494 5128 81154 352840
rect 81934 5128 84874 352840
rect 85654 5128 88594 352840
rect 89374 5128 96034 352840
rect 96814 5128 99754 352840
rect 100534 5128 109714 352840
rect 110494 5128 113434 352840
rect 114214 5128 117154 352840
rect 117934 5128 120874 352840
rect 121654 5128 124594 352840
rect 125374 5128 128314 352840
rect 129094 5128 132034 352840
rect 132814 5128 135754 352840
rect 136534 5128 145714 352840
rect 146494 5128 149434 352840
rect 150214 5128 153154 352840
rect 153934 5128 156874 352840
rect 157654 5128 160594 352840
rect 161374 5128 164314 352840
rect 165094 5128 168034 352840
rect 168814 5128 171754 352840
rect 172534 5128 181714 352840
rect 182494 5128 189154 352840
rect 189934 5128 192874 352840
rect 193654 5128 196594 352840
rect 197374 5128 204034 352840
rect 204814 5128 207754 352840
rect 208534 5128 217714 352840
rect 218494 5128 221434 352840
rect 222214 5128 225154 352840
rect 225934 5128 228874 352840
rect 229654 5128 232594 352840
rect 233374 5128 236314 352840
rect 237094 5128 240034 352840
rect 240814 5128 243754 352840
rect 244534 5128 253714 352840
rect 254494 5128 257434 352840
rect 258214 5128 264874 352840
rect 265654 5128 268594 352840
rect 269374 5128 272314 352840
rect 273094 5128 276034 352840
rect 276814 5128 279754 352840
rect 280534 5128 289714 352840
rect 290494 5128 293434 352840
rect 294214 5128 297154 352840
rect 297934 5128 300874 352840
rect 301654 5128 304594 352840
rect 305374 5128 312034 352840
rect 312814 5128 315754 352840
rect 316534 5128 325714 352840
rect 326494 5128 329434 352840
rect 330214 5128 333154 352840
rect 333934 5128 336874 352840
rect 337654 5128 340594 352840
rect 341374 5128 344314 352840
rect 345094 5128 348034 352840
rect 348814 5128 351754 352840
rect 352534 5128 361714 352840
rect 362494 5128 365434 352840
rect 366214 5128 372874 352840
rect 373654 5128 376594 352840
rect 377374 5128 380314 352840
rect 381094 5128 387754 352840
rect 388534 5128 397714 352840
rect 398494 5128 401434 352840
rect 402214 5128 405154 352840
rect 405934 5128 408874 352840
rect 409654 5128 412594 352840
rect 413374 5128 416314 352840
rect 417094 5128 420034 352840
rect 420814 5128 423754 352840
rect 424534 5128 433714 352840
rect 434494 5128 437434 352840
rect 438214 5128 441154 352840
rect 441934 5128 444874 352840
rect 445654 5128 448594 352840
rect 449374 5128 452314 352840
rect 453094 5128 456034 352840
rect 456814 5128 459754 352840
rect 460534 5128 469714 352840
rect 470494 5128 473434 352840
rect 474214 5128 480874 352840
rect 481654 5128 484594 352840
rect 485374 5128 488314 352840
rect 489094 5128 495754 352840
rect 496534 5128 505714 352840
rect 506494 5128 509434 352840
rect 510214 5128 513154 352840
rect 513934 5128 516874 352840
rect 517654 5128 520594 352840
rect 521374 5128 524314 352840
rect 525094 5128 528034 352840
rect 528814 5128 531754 352840
rect 532534 5128 541714 352840
rect 542494 5128 545434 352840
rect 546214 5128 549154 352840
rect 549934 5128 552874 352840
rect 553654 5128 556594 352840
rect 557374 5128 560314 352840
rect 561094 5128 564034 352840
rect 564814 5128 567754 352840
rect 568534 5128 569488 352840
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 698026 592650 698646
rect -8726 694306 592650 694926
rect -8726 690586 592650 691206
rect -8726 686866 592650 687486
rect -8726 676906 592650 677526
rect -8726 673186 592650 673806
rect -8726 669466 592650 670086
rect -8726 665746 592650 666366
rect -8726 662026 592650 662646
rect -8726 658306 592650 658926
rect -8726 654586 592650 655206
rect -8726 650866 592650 651486
rect -8726 640906 592650 641526
rect -8726 637186 592650 637806
rect -8726 633466 592650 634086
rect -8726 629746 592650 630366
rect -8726 626026 592650 626646
rect -8726 622306 592650 622926
rect -8726 618586 592650 619206
rect -8726 614866 592650 615486
rect -8726 604906 592650 605526
rect -8726 601186 592650 601806
rect -8726 597466 592650 598086
rect -8726 593746 592650 594366
rect -8726 590026 592650 590646
rect -8726 586306 592650 586926
rect -8726 582586 592650 583206
rect -8726 578866 592650 579486
rect -8726 568906 592650 569526
rect -8726 565186 592650 565806
rect -8726 561466 592650 562086
rect -8726 557746 592650 558366
rect -8726 554026 592650 554646
rect -8726 550306 592650 550926
rect -8726 546586 592650 547206
rect -8726 542866 592650 543486
rect -8726 532906 592650 533526
rect -8726 529186 592650 529806
rect -8726 525466 592650 526086
rect -8726 521746 592650 522366
rect -8726 518026 592650 518646
rect -8726 514306 592650 514926
rect -8726 510586 592650 511206
rect -8726 506866 592650 507486
rect -8726 496906 592650 497526
rect -8726 493186 592650 493806
rect -8726 489466 592650 490086
rect -8726 485746 592650 486366
rect -8726 482026 592650 482646
rect -8726 478306 592650 478926
rect -8726 474586 592650 475206
rect -8726 470866 592650 471486
rect -8726 460906 592650 461526
rect -8726 457186 592650 457806
rect -8726 453466 592650 454086
rect -8726 449746 592650 450366
rect -8726 446026 592650 446646
rect -8726 442306 592650 442926
rect -8726 438586 592650 439206
rect -8726 434866 592650 435486
rect -8726 424906 592650 425526
rect -8726 421186 592650 421806
rect -8726 417466 592650 418086
rect -8726 413746 592650 414366
rect -8726 410026 592650 410646
rect -8726 406306 592650 406926
rect -8726 402586 592650 403206
rect -8726 398866 592650 399486
rect -8726 388906 592650 389526
rect -8726 385186 592650 385806
rect -8726 381466 592650 382086
rect -8726 377746 592650 378366
rect -8726 374026 592650 374646
rect -8726 370306 592650 370926
rect -8726 366586 592650 367206
rect -8726 362866 592650 363486
rect -8726 352906 592650 353526
rect -8726 349186 592650 349806
rect -8726 345466 592650 346086
rect -8726 341746 592650 342366
rect -8726 338026 592650 338646
rect -8726 334306 592650 334926
rect -8726 330586 592650 331206
rect -8726 326866 592650 327486
rect -8726 316906 592650 317526
rect -8726 313186 592650 313806
rect -8726 309466 592650 310086
rect -8726 305746 592650 306366
rect -8726 302026 592650 302646
rect -8726 298306 592650 298926
rect -8726 294586 592650 295206
rect -8726 290866 592650 291486
rect -8726 280906 592650 281526
rect -8726 277186 592650 277806
rect -8726 273466 592650 274086
rect -8726 269746 592650 270366
rect -8726 266026 592650 266646
rect -8726 262306 592650 262926
rect -8726 258586 592650 259206
rect -8726 254866 592650 255486
rect -8726 244906 592650 245526
rect -8726 241186 592650 241806
rect -8726 237466 592650 238086
rect -8726 233746 592650 234366
rect -8726 230026 592650 230646
rect -8726 226306 592650 226926
rect -8726 222586 592650 223206
rect -8726 218866 592650 219486
rect -8726 208906 592650 209526
rect -8726 205186 592650 205806
rect -8726 201466 592650 202086
rect -8726 197746 592650 198366
rect -8726 194026 592650 194646
rect -8726 190306 592650 190926
rect -8726 186586 592650 187206
rect -8726 182866 592650 183486
rect -8726 172906 592650 173526
rect -8726 169186 592650 169806
rect -8726 165466 592650 166086
rect -8726 161746 592650 162366
rect -8726 158026 592650 158646
rect -8726 154306 592650 154926
rect -8726 150586 592650 151206
rect -8726 146866 592650 147486
rect -8726 136906 592650 137526
rect -8726 133186 592650 133806
rect -8726 129466 592650 130086
rect -8726 125746 592650 126366
rect -8726 122026 592650 122646
rect -8726 118306 592650 118926
rect -8726 114586 592650 115206
rect -8726 110866 592650 111486
rect -8726 100906 592650 101526
rect -8726 97186 592650 97806
rect -8726 93466 592650 94086
rect -8726 89746 592650 90366
rect -8726 86026 592650 86646
rect -8726 82306 592650 82926
rect -8726 78586 592650 79206
rect -8726 74866 592650 75486
rect -8726 64906 592650 65526
rect -8726 61186 592650 61806
rect -8726 57466 592650 58086
rect -8726 53746 592650 54366
rect -8726 50026 592650 50646
rect -8726 46306 592650 46926
rect -8726 42586 592650 43206
rect -8726 38866 592650 39486
rect -8726 28906 592650 29526
rect -8726 25186 592650 25806
rect -8726 21466 592650 22086
rect -8726 17746 592650 18366
rect -8726 14026 592650 14646
rect -8726 10306 592650 10926
rect -8726 6586 592650 7206
rect -8726 2866 592650 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 1 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 2 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 3 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 4 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 5 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 6 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 7 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 8 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 9 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 10 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 11 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 12 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 13 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 14 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 15 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 16 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 17 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 18 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 19 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 20 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 21 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 22 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 23 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 24 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 25 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 26 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 27 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 28 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 29 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 30 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 31 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 32 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 33 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 34 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 35 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 36 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 37 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 38 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 39 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 40 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 41 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 42 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 43 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 44 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 45 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 46 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 47 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 48 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 49 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 50 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 51 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 52 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 53 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 54 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 55 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 56 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 57 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 58 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 59 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 60 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 61 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 62 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 63 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 64 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 65 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 66 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 67 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 68 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 69 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 70 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 71 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 72 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 73 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 74 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 75 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 76 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 77 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 78 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 79 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 80 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 81 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 82 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 83 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 84 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 85 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 86 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 87 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 88 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 89 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 90 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 91 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 92 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 93 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 94 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 95 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 96 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 97 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 98 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 99 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 100 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 101 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 102 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 103 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 104 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 105 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 106 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 107 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 108 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 109 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 110 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 111 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 112 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 113 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 114 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 115 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 116 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 117 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 118 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 119 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 120 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 121 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 122 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 123 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 124 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 125 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 126 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 127 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 128 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 129 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 130 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 131 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 132 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 133 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 134 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 135 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 136 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 137 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 138 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 139 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 140 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 141 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 142 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 143 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 144 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 145 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 146 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 147 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 148 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 149 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 150 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 151 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 152 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 153 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 154 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 155 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 156 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 157 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 158 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 159 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 160 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 161 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 162 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 163 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 164 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 165 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 166 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 167 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 168 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 169 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 170 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 171 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 172 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 173 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 174 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 175 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 176 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 177 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 178 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 179 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 180 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 181 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 182 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 183 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 184 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 185 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 186 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 187 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 188 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 189 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 190 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 191 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 192 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 193 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 194 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 195 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 196 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 197 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 198 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 199 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 200 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 201 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 202 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 203 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 204 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 205 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 206 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 207 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 208 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 209 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 210 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 211 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 212 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 213 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 214 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 215 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 216 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 217 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 218 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 219 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 220 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 221 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 222 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 223 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 224 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 225 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 226 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 227 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 228 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 229 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 230 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 231 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 232 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 233 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 234 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 235 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 236 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 237 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 238 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 239 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 240 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 241 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 242 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 243 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 244 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 245 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 246 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 247 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 248 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 249 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 250 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 251 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 252 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 253 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 254 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 255 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 256 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 257 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 257 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 9234 -7654 9854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 45234 -7654 45854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 81234 -7654 81854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 117234 -7654 117854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 153234 -7654 153854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 189234 -7654 189854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 225234 -7654 225854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 261234 354980 261854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 297234 -7654 297854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 333234 -7654 333854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 369234 354980 369854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 405234 -7654 405854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 441234 -7654 441854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 477234 354980 477854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 513234 -7654 513854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s 549234 -7654 549854 711590 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 10306 592650 10926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 46306 592650 46926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 82306 592650 82926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 118306 592650 118926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 154306 592650 154926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 190306 592650 190926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 226306 592650 226926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 262306 592650 262926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 298306 592650 298926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 334306 592650 334926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 370306 592650 370926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 406306 592650 406926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 442306 592650 442926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 478306 592650 478926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 514306 592650 514926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 550306 592650 550926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 586306 592650 586926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 622306 592650 622926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 658306 592650 658926 6 vccd2
port 258 nsew power bidirectional
rlabel metal5 s -8726 694306 592650 694926 6 vccd2
port 258 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 16674 -7654 17294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 52674 -7654 53294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 88674 -7654 89294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 124674 -7654 125294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 160674 -7654 161294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 196674 -7654 197294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 232674 -7654 233294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 268674 -7654 269294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 304674 -7654 305294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 340674 -7654 341294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 376674 -7654 377294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 412674 -7654 413294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 448674 -7654 449294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 484674 -7654 485294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 520674 -7654 521294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s 556674 -7654 557294 711590 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 17746 592650 18366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 53746 592650 54366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 89746 592650 90366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 125746 592650 126366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 161746 592650 162366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 197746 592650 198366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 233746 592650 234366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 269746 592650 270366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 305746 592650 306366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 341746 592650 342366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 377746 592650 378366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 413746 592650 414366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 449746 592650 450366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 485746 592650 486366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 521746 592650 522366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 557746 592650 558366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 593746 592650 594366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 629746 592650 630366 6 vdda1
port 259 nsew power bidirectional
rlabel metal5 s -8726 665746 592650 666366 6 vdda1
port 259 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 24114 -7654 24734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 60114 -7654 60734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 96114 -7654 96734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 132114 -7654 132734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 168114 -7654 168734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 204114 -7654 204734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 240114 -7654 240734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 276114 -7654 276734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 312114 -7654 312734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 348114 -7654 348734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 384114 354980 384734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 420114 -7654 420734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 456114 -7654 456734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 492114 354980 492734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 528114 -7654 528734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 564114 -7654 564734 711590 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 25186 592650 25806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 61186 592650 61806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 97186 592650 97806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 133186 592650 133806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 169186 592650 169806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 205186 592650 205806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 241186 592650 241806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 277186 592650 277806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 313186 592650 313806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 349186 592650 349806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 385186 592650 385806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 421186 592650 421806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 457186 592650 457806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 493186 592650 493806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 529186 592650 529806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 565186 592650 565806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 601186 592650 601806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 637186 592650 637806 6 vdda2
port 260 nsew power bidirectional
rlabel metal5 s -8726 673186 592650 673806 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 20394 -7654 21014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 56394 -7654 57014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 92394 354980 93014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 128394 -7654 129014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 164394 -7654 165014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 200394 354980 201014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 236394 -7654 237014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 272394 -7654 273014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 308394 354980 309014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 344394 -7654 345014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 380394 -7654 381014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 416394 -7654 417014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 452394 -7654 453014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 488394 -7654 489014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 524394 -7654 525014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 560394 -7654 561014 711590 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 21466 592650 22086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 57466 592650 58086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 93466 592650 94086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 129466 592650 130086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 165466 592650 166086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 201466 592650 202086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 237466 592650 238086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 273466 592650 274086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 309466 592650 310086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 345466 592650 346086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 381466 592650 382086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 417466 592650 418086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 453466 592650 454086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 489466 592650 490086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 525466 592650 526086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 561466 592650 562086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 597466 592650 598086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 633466 592650 634086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal5 s -8726 669466 592650 670086 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 27834 -7654 28454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 63834 -7654 64454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 99834 -7654 100454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 135834 -7654 136454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 171834 -7654 172454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 207834 -7654 208454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 243834 -7654 244454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 279834 -7654 280454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 315834 -7654 316454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 351834 -7654 352454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 387834 -7654 388454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 423834 -7654 424454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 459834 -7654 460454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 495834 -7654 496454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 531834 -7654 532454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s 567834 -7654 568454 711590 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 28906 592650 29526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 64906 592650 65526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 100906 592650 101526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 136906 592650 137526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 172906 592650 173526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 208906 592650 209526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 244906 592650 245526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 280906 592650 281526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 316906 592650 317526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 352906 592650 353526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 388906 592650 389526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 424906 592650 425526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 460906 592650 461526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 496906 592650 497526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 532906 592650 533526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 568906 592650 569526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 604906 592650 605526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 640906 592650 641526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal5 s -8726 676906 592650 677526 6 vssa2
port 262 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 5514 -7654 6134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 41514 -7654 42134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 77514 354980 78134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 113514 -7654 114134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 149514 -7654 150134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 185514 354980 186134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 221514 -7654 222134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 257514 -7654 258134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 293514 -7654 294134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 329514 -7654 330134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 365514 -7654 366134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 401514 -7654 402134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 437514 -7654 438134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 473514 -7654 474134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 509514 -7654 510134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 545514 -7654 546134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 581514 -7654 582134 711590 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 6586 592650 7206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 42586 592650 43206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 78586 592650 79206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 114586 592650 115206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 150586 592650 151206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 186586 592650 187206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 222586 592650 223206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 258586 592650 259206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 294586 592650 295206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 330586 592650 331206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 366586 592650 367206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 402586 592650 403206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 438586 592650 439206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 474586 592650 475206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 510586 592650 511206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 546586 592650 547206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 582586 592650 583206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 618586 592650 619206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 654586 592650 655206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -8726 690586 592650 691206 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 12954 -7654 13574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 48954 -7654 49574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 84954 -7654 85574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 120954 -7654 121574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 156954 -7654 157574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 192954 -7654 193574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 228954 -7654 229574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 264954 -7654 265574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 300954 -7654 301574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 336954 -7654 337574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 372954 -7654 373574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 408954 -7654 409574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 444954 -7654 445574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 480954 -7654 481574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 516954 -7654 517574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal4 s 552954 -7654 553574 711590 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 14026 592650 14646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 50026 592650 50646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 86026 592650 86646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 122026 592650 122646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 158026 592650 158646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 194026 592650 194646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 230026 592650 230646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 266026 592650 266646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 302026 592650 302646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 338026 592650 338646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 374026 592650 374646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 410026 592650 410646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 446026 592650 446646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 482026 592650 482646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 518026 592650 518646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 554026 592650 554646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 590026 592650 590646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 626026 592650 626646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 662026 592650 662646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal5 s -8726 698026 592650 698646 6 vssd2
port 264 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 265 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 266 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 52634518
string GDS_FILE /home/vboxuser/Documents/samj_user_project/openlane/user_project_wrapper/runs/24_10_23_21_55/results/signoff/user_project_wrapper.magic.gds
string GDS_START 51502396
<< end >>

